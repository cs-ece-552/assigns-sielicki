module DataMemory {

}
