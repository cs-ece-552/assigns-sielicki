module xnor5_1(
  input  [4:0] func,
  input  [4:0] opcode,
  output       out
);
  wire  _GEN_0;
  wire  _GEN_1;
  wire  _GEN_2;
  wire  _xor_____verilog_xnor5_1_v_7_1027;
  wire  xor0;
  wire  _GEN_3;
  wire  _GEN_4;
  wire  _GEN_5;
  wire  _xor_____verilog_xnor5_1_v_8_1029;
  wire  xor1;
  wire  _GEN_6;
  wire  _and_____verilog_xnor5_1_v_13_1037;
  wire  _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire  _xor_____verilog_xnor5_1_v_9_1031;
  wire  xor2;
  wire  _GEN_10;
  wire  _and_____verilog_xnor5_1_v_13_1038;
  wire  _GEN_11;
  wire  _GEN_12;
  wire  _GEN_13;
  wire  _xor_____verilog_xnor5_1_v_10_1033;
  wire  xor3;
  wire  _GEN_14;
  wire  _and_____verilog_xnor5_1_v_13_1039;
  wire  _GEN_15;
  wire  _GEN_16;
  wire  _GEN_17;
  wire  _xor_____verilog_xnor5_1_v_11_1035;
  wire  xor4;
  wire  _GEN_18;
  assign _GEN_0 = func[0];
  assign _GEN_1 = opcode[0];
  assign _GEN_2 = $unsigned(_GEN_0);
  assign _xor_____verilog_xnor5_1_v_7_1027 = _GEN_1 ^ _GEN_2;
  assign xor0 = ~ _xor_____verilog_xnor5_1_v_7_1027;
  assign _GEN_3 = func[1];
  assign _GEN_4 = opcode[1];
  assign _GEN_5 = $unsigned(_GEN_3);
  assign _xor_____verilog_xnor5_1_v_8_1029 = _GEN_4 ^ _GEN_5;
  assign xor1 = ~ _xor_____verilog_xnor5_1_v_8_1029;
  assign _GEN_6 = $unsigned(xor1);
  assign _and_____verilog_xnor5_1_v_13_1037 = xor0 & _GEN_6;
  assign _GEN_7 = func[2];
  assign _GEN_8 = opcode[2];
  assign _GEN_9 = $unsigned(_GEN_7);
  assign _xor_____verilog_xnor5_1_v_9_1031 = _GEN_8 ^ _GEN_9;
  assign xor2 = ~ _xor_____verilog_xnor5_1_v_9_1031;
  assign _GEN_10 = $unsigned(xor2);
  assign _and_____verilog_xnor5_1_v_13_1038 = _and_____verilog_xnor5_1_v_13_1037 & _GEN_10;
  assign _GEN_11 = func[3];
  assign _GEN_12 = opcode[3];
  assign _GEN_13 = $unsigned(_GEN_11);
  assign _xor_____verilog_xnor5_1_v_10_1033 = _GEN_12 ^ _GEN_13;
  assign xor3 = ~ _xor_____verilog_xnor5_1_v_10_1033;
  assign _GEN_14 = $unsigned(xor3);
  assign _and_____verilog_xnor5_1_v_13_1039 = _and_____verilog_xnor5_1_v_13_1038 & _GEN_14;
  assign _GEN_15 = func[4];
  assign _GEN_16 = opcode[4];
  assign _GEN_17 = $unsigned(_GEN_15);
  assign _xor_____verilog_xnor5_1_v_11_1035 = _GEN_16 ^ _GEN_17;
  assign xor4 = ~ _xor_____verilog_xnor5_1_v_11_1035;
  assign _GEN_18 = $unsigned(xor4);
  assign out = _and_____verilog_xnor5_1_v_13_1039 & _GEN_18;
endmodule
